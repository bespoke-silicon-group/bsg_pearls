
// replace with hardened buffer with decent drive strength
module bsg_clk_gen_monitor_clk_buf
  (input          i
   , output logic o
   );

  assign o = i;

endmodule

